* ��Ŀ D:\work\pads\gps\sch\gps.cir
* ���� Mentor Graphics ��·���汾 1.0.0
* Inifile   : 
* Options   : 

* ����Ԫ���� C1 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C2 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C3 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C4 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C5 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C6 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C7 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�
* ����Ԫ���� C8 ������Ϊδ�ҵ� Sim.Analog.Prefix ���ԡ�

.END
